module my_xor(
  input a,
  input b,
  output out
  );
  xor w1(out,a,b);
  
endmodule