module ALU_test;
reg signed [63:0] a,b;
reg [1:0] mg_op;
wire signed [63:0] c;
wire overflow;

ALU A1 (overflow,c,a,b, mg_op);
initial
begin
  $dumpfile("ALU_gtk.vcd");
  $dumpvars;
   a = 64'b111111111111111111111111110000111111111111111111111111111111; b=64'b111111111111000011111111111111111111111111111111111111111111; mg_op= 2'b00;
  #5 a = 64'b011111111111111111111111111111111111111100001111111111111111; b=64'b011111111111111111111111111111111111111111111100001111111111;  mg_op = 2'b01;
  #5 a = 64'b011111111111111111000011111111111111111111111111111111111111; b=64'b111111111111111111111111111111111000011111111111111111111111;  mg_op = 2'b10;
  #5 a = 64'b100000000000000000000000000000000000000000000000000000000001; b=64'b1111111111111111100001111111111111111111111111111111111111100000;mg_op = 2'b11;
  #10 $finish;
end

initial begin
$display ("Control = 0 --> ADD");  
$display ("Control = 1 --> SUB");  
$display ("Control = 2 --> AND");  
$display ("Control = 3 --> XOR\n");  
end

initial 
	$monitor("Control = %d\n a  = %d\n b  = %d\noverflow = %b\n c  = %d\n",mg_op,a,b,overflow,c);
endmodule

