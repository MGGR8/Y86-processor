module my_and(
  input a,
  input b,
  output out
  );
  and w1(out,a,b);
  
endmodule